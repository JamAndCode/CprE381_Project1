-------------------------------------------------------------------------
-- Jamie Anderson
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- 5to32_decode.vhd
----------------------------------------------------------------------------
-- DESCRIPTION: This file contains a 5-to-32 bit decoder for a MIPS register
----------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

entity decode_5to32 is
  port( i_Enable: in std_logic;
	i_A	: in std_logic_vector(4 downto 0);
	o_F	: out std_logic_vector(31 downto 0));
end decode_5to32;

architecture dataflow of decode_5to32 is
begin

	process(i_Enable, i_A) is
	begin
	if (i_Enable = '1') then
	case i_A is
		when  "00000" => o_F <= "00000000000000000000000000000001";
		when  "00001" => o_F <=  "00000000000000000000000000000010";
		when  "00010" => o_F <= "00000000000000000000000000000100";
		when  "00011" => o_F <= "00000000000000000000000000001000";
		when  "00100" => o_F <= "00000000000000000000000000010000";
		when  "00101" => o_F <=  "00000000000000000000000000100000";
		when  "00110" => o_F <= "00000000000000000000000001000000";
		when  "00111" => o_F <= "00000000000000000000000010000000";
		when "01000" => o_F <= "00000000000000000000000100000000" ;
		when "01001" => o_F <= "00000000000000000000001000000000";
		when "01010" => o_F <= "00000000000000000000010000000000";
		when  "01011" => o_F <= "00000000000000000000100000000000";
		when  "01100" => o_F <= "00000000000000000001000000000000";
		when  "01101" => o_F <= "00000000000000000010000000000000";
		when  "01110" => o_F <=  "00000000000000000100000000000000";
		when  "01111" => o_F <= "00000000000000001000000000000000";
		when  "10000" => o_F <= "00000000000000010000000000000000";
		when  "10001" => o_F <= "00000000000000100000000000000000";
		when  "10010" => o_F <= "00000000000001000000000000000000";
		when  "10011" => o_F <= "00000000000010000000000000000000";
		when  "10100" => o_F <= "00000000000100000000000000000000";
		when  "10101" => o_F <=  "00000000001000000000000000000000";
		when  "10110" => o_F <=  "00000000010000000000000000000000";
		when  "10111" => o_F <=  "00000000100000000000000000000000";
		when  "11000" => o_F <=  "00000001000000000000000000000000";
		when  "11001" => o_F <=  "00000010000000000000000000000000";
		when  "11010" => o_F <= "00000100000000000000000000000000" ;
		when  "11011" => o_F <=  "00001000000000000000000000000000";
		when  "11100" => o_F <= "00010000000000000000000000000000";
		when  "11101" => o_F <= "00100000000000000000000000000000";
		when  "11110" => o_F <= "01000000000000000000000000000000";
		when  "11111" => o_F <= "10000000000000000000000000000000";
		when others => o_F <=  "00000000000000000000000000000000";
		end case;
		else
			o_F <= "00000000000000000000000000000000";
end if;
	end process;
end dataflow;
